* C:\Users\lenovo\eSim-Workspace\sinewave_generator\sinewave_generator.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 03/17/21 16:41:33

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  Net-_U1-Pad1_ ? in Net-_U1-Pad4_ dff		
U2  Net-_U1-Pad4_ ? in Net-_U2-Pad4_ dff		
U5  Net-_U2-Pad4_ ? in Net-_U5-Pad4_ dff		
U6  Net-_U5-Pad4_ ? in Net-_U6-Pad4_ dff		
U9  Net-_U6-Pad4_ Net-_U1-Pad1_ d_inverter		
U4  Net-_U4-Pad1_ in adc_bridge_1		
U7  Net-_U1-Pad4_ Net-_U2-Pad4_ Net-_U5-Pad4_ Net-_R1-Pad2_ Net-_R2-Pad2_ Net-_R3-Pad2_ dac_bridge_3		
R1  out Net-_R1-Pad2_ 10k		
R2  out Net-_R2-Pad2_ 20k		
R3  out Net-_R3-Pad2_ 10k		
U8  out plot_v1		
U3  in plot_v1		
v1  Net-_U4-Pad1_ GND 5v		

.end
